LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE ieee.std_logic_textio.ALL;
USE std.textio.ALL;

ENTITY Memory IS
    GENERIC (
        DATA_WIDTH : INTEGER := 32;
        ADDR_WIDTH : INTEGER := 10; -- 1024 memory locations
        INIT_FILE : STRING := ""
    );
    PORT (
        clk : IN STD_LOGIC;
        write_enable : IN STD_LOGIC;
        address : IN STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);
        data_in : IN STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
        data_out : OUT STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0)
    );
END Memory;

ARCHITECTURE Beh OF Memory IS
    TYPE memory_array IS ARRAY (0 TO (2 ** ADDR_WIDTH) - 1) OF STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
    -- PY_START_EDITING
    SIGNAL memory : memory_array := (
    0 => "00000100000000010000000000000101", -- LI R1, 5
    1 => "00000100000000100000000000000110", -- LI R2, 6
    2 => "00000000001000100001100000000010", -- ADD R3, R1, R2
    3 => "00001000000000110000000000000000", -- OUT R3
    4 => "00000100000001000000000000000111", -- LI R4, 7
    5 => "00000000001001000010100000000001", -- XOR R5, R1, R4
    6 => "00001000000001010000000000000000", -- OUT R5
    7 => "00000000000000010011000010000110", -- LSL R6, R1, 2
    8 => "00001000000001100000000000000000", -- OUT R6
    9 => "00000100000000100000000000010000", -- LI R2, 16
    10 => "00000000000000100011100010000111", -- LSR R7, R2, 2
    11 => "00001000000001110000000000000000", -- OUT R7
    OTHERS => (OTHERS => '0')
    );
    -- PY_END_EDITING

BEGIN
    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            IF write_enable = '1' THEN
                memory(to_integer(unsigned(address))) <= data_in;
            END IF;
        END IF;
    END PROCESS;
    data_out <= memory(to_integer(unsigned(address)));
END ARCHITECTURE;